`timescale 1ns / 1ps
//Master controller
 module ctrl(e,op,funct,RegWrite,ALUSrc,RegDst,MemtoReg,MemWrite,NPCCtrl,ExtOp,aluc,MA3D,MALUOUT);
input[5:0] op,funct;
input e;
output[1:0] NPCCtrl;
output[2:0] aluc;
output RegWrite,ALUSrc,RegDst,MemtoReg,ExtOp,MemWrite,MA3D,MALUOUT;

reg[1:0] NPCCtrl=0;
reg[2:0] aluc=0;
reg RegWrite=0,ALUSrc=0,RegDst=0,MemtoReg=0,ExtOp=0,MemWrite=0,MA3D=0,MALUOUT=0;

always @ (e,op,funct)
begin
   if(e==1)//stall
	begin
	   RegWrite<=0;
		ALUSrc<=0;
		RegDst<=0;
		MemtoReg<=0;
		MemWrite<=0;
		NPCCtrl<=2'b00;
		ExtOp<=0;
		aluc<=3'b000;
		MA3D<=0;
		MALUOUT<=0;
	end
	else
	begin
		case(op)
		/*6'b001110://XORI
		begin
			RegWrite<=1;
			ALUSrc<=1;
			RegDst<=0;
			MemtoReg<=0;
			MemWrite<=0;
			NPCCtrl<=2'b00;
			ExtOp<=0;
			aluc<=3'b011;
			MA3D<=0;
		end*/
		6'b000000:
		begin	
			ALUSrc<=0;
			RegDst<=1;
			MemtoReg<=0;
			MemWrite<=0;
			ExtOp<=0;
			MA3D<=0;
			MALUOUT<=0;
			case(funct)
			6'b100001://ADDU
			begin
				NPCCtrl<=2'b00;
				RegWrite<=1;
				aluc<=3'b010;
			end
			6'b000000://NOP
			begin
				NPCCtrl<=2'b00;
				RegWrite<=0;
				aluc<=3'b100;
			end
			6'b001000://JR
			begin
				NPCCtrl<=2'b11;
				RegWrite<=0;
				aluc<=3'b111;
			end
			6'b100011://SUBU
			begin
				NPCCtrl<=2'b00;
				RegWrite<=1;
				aluc<=3'b110;
			end
			6'b100100://AND
			begin
				NPCCtrl<=2'b00;
				RegWrite<=1;
				aluc<=3'b000;
			end
			6'b100101://OR
			begin
				NPCCtrl<=2'b00;
				RegWrite<=1;
				aluc<=3'b001;
			end
			endcase
		end
		6'b001101://ORI
		begin
			RegWrite<=1;
			ALUSrc<=1;
			RegDst<=0;
			MemtoReg<=0;
			MemWrite<=0;
			NPCCtrl<=2'b00;
			ExtOp<=0;
			aluc<=3'b001;
			MA3D<=0;
			MALUOUT<=0;
		end
		6'b100011://LW
		begin
			RegWrite<=1;
			ALUSrc<=1;
			RegDst<=0;
			MemtoReg<=1;
			MemWrite<=0;
			NPCCtrl<=2'b00;
			ExtOp<=1;
			aluc<=3'b010;
			MA3D<=0;
			MALUOUT<=0;
		end
		6'b101011://SW
		begin
			RegWrite<=0;
			ALUSrc<=1;
			RegDst<=0;
			MemtoReg<=0;
			MemWrite<=1;
			NPCCtrl<=2'b00;
			ExtOp<=1;
			aluc<=3'b010;
			MA3D<=0;
			MALUOUT<=0;
		end
		6'b000100://BEQ
		begin
			RegWrite<=0;
			ALUSrc<=0;
			RegDst<=0;
			MemtoReg<=0;
			MemWrite<=0;
			NPCCtrl<=2'b10;
			ExtOp<=0;
			aluc<=3'b111;
			MA3D<=0;
			MALUOUT<=0;
		end
		6'b000010://J
		begin
			RegWrite<=0;
			ALUSrc<=0;
			RegDst<=0;
			MemtoReg<=0;
			MemWrite<=0;
			NPCCtrl<=2'b01;
			ExtOp<=0;
			aluc<=3'b111;
			MA3D<=0;
			MALUOUT<=0;
		end
		6'b000011://JAL
		begin
			RegWrite<=1;
			ALUSrc<=0;
			RegDst<=0;
			MemtoReg<=0;
			MemWrite<=0;
			NPCCtrl<=2'b01;
			ExtOp<=0;
			aluc<=3'b111;
			MA3D<=1;
			MALUOUT<=1;
		end
		6'b001111://LUI
		begin
			RegWrite<=1;
			ALUSrc<=1;
			RegDst<=0;
			MemtoReg<=0;
			MemWrite<=0;
			NPCCtrl<=2'b00;
			ExtOp<=0;
			aluc<=3'b100;
			MA3D<=0;
			MALUOUT<=0;
		end
		6'b001000://ADDI
		begin
			RegWrite<=1;
			ALUSrc<=1;
			RegDst<=0;
			MemtoReg<=0;
			MemWrite<=0;
			NPCCtrl<=2'b00;
			ExtOp<=0;
			aluc<=3'b010;
			MA3D<=0;
			MALUOUT<=0;
		end
		endcase
	end
end

endmodule
